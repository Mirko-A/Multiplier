----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/14/2021 09:33:01 PM
-- Design Name: 
-- Module Name: pipo_reg - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pipo_reg is
    generic (WIDTH: positive := 8);
    Port ( d : in STD_LOGIC_VECTOR(WIDTH-1 downto 0);
           clk : in STD_LOGIC;
           q : out STD_LOGIC_VECTOR(WIDTH-1 downto 0));
end pipo_reg;

architecture Behavioral of pipo_reg is

begin
    
    reg: process (clk) is 
        begin
            if(clk'event and clk='1') then
                q <= d;
            end if;
        end process;

end Behavioral;
